library verilog;
use verilog.vl_types.all;
entity cont_productos_vlg_vec_tst is
end cont_productos_vlg_vec_tst;
