library verilog;
use verilog.vl_types.all;
entity capacidad_val_vlg_check_tst is
    port(
        capacidad       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end capacidad_val_vlg_check_tst;
