library verilog;
use verilog.vl_types.all;
entity digitos_vlg_vec_tst is
end digitos_vlg_vec_tst;
