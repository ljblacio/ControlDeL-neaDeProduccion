library verilog;
use verilog.vl_types.all;
entity valor_pwm_vlg_vec_tst is
end valor_pwm_vlg_vec_tst;
