library verilog;
use verilog.vl_types.all;
entity frec_var_vlg_check_tst is
    port(
        frec            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end frec_var_vlg_check_tst;
