library verilog;
use verilog.vl_types.all;
entity separa_3dig_vlg_vec_tst is
end separa_3dig_vlg_vec_tst;
