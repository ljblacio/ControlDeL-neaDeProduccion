library verilog;
use verilog.vl_types.all;
entity separador_3dig_vlg_vec_tst is
end separador_3dig_vlg_vec_tst;
