library verilog;
use verilog.vl_types.all;
entity capacidad_val_vlg_vec_tst is
end capacidad_val_vlg_vec_tst;
