library verilog;
use verilog.vl_types.all;
entity CONTROL_PRODUCCION_SIMULAR_vlg_vec_tst is
end CONTROL_PRODUCCION_SIMULAR_vlg_vec_tst;
