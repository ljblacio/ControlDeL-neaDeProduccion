library verilog;
use verilog.vl_types.all;
entity frec_var_vlg_vec_tst is
end frec_var_vlg_vec_tst;
