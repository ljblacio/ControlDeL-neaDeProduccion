library verilog;
use verilog.vl_types.all;
entity cont_updw_vlg_vec_tst is
end cont_updw_vlg_vec_tst;
